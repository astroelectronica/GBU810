.title KiCad schematic
.include "C:/AE/GBU810/_models/GBU810.spice.txt"
C1 /VBULK 0 {CBULK}
I1 /VOUT 0 {ILOAD}
R1 /VOUT /VBULK {RSER}
D3 0 /LINE DI_GBU810
D4 0 /NEUTRAL DI_GBU810
D2 /NEUTRAL /VOUT DI_GBU810
D1 /LINE /VOUT DI_GBU810
V1 /LINE /NEUTRAL SINE({VOFFSET} {VPK} {FREQ})
.end
